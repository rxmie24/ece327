library ieee;
use ieee.std_logic_1164.all;

-- insert entity definition here

-- insert architecture here

-- test comment

